parameter WIDTH = 32;
parameter DEPTH = 4;
